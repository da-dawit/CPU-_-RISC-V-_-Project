module rf (
    input              clk,
    input              we,
    input      [4:0]   rs1,
    input      [4:0]   rs2,
    input      [4:0]   rd,
    input      [31:0]  wd,
    output     [31:0]  rd1,
    output     [31:0]  rd2
);

    reg [31:0] regs [31:0];
    
    // Initialize all registers to 0
    integer i;
    initial begin
        for (i = 0; i < 32; i = i + 1)
            regs[i] = 32'h00000000;
    end

    // READ PORTS: combinational
    assign rd1 = (rs1 == 0) ? 32'b0 : regs[rs1];
    assign rd2 = (rs2 == 0) ? 32'b0 : regs[rs2];

    // WRITE PORT: synchronous
    always @(posedge clk) begin
        if (we && (rd != 0))
            regs[rd] <= wd;
    end

endmodule